/* Linda Zhang
    AHB access point with connection to generic bus design 
*/ 

`include "ahb_ap_if.vh"
`include "jtag_types_pkg.vh"

module ahb_ap_generic_bus (
    
);
    
endmodule