/* Wen-Bo Hung, created at 2023/11/2, email: hong395@purdue.edu, peterhouse08271026@gmail.com*/
// JTAG SoCET Team
// Instruction decoder

